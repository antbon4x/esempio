version https://git-lfs.github.com/spec/v1
oid sha256:52081b4cb0ee6236a12e8a9116a23fd6811277a47619f90cc8224d442a071898
size 6757
