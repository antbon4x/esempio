version https://git-lfs.github.com/spec/v1
oid sha256:7d3b73b91faafeb483a306ea5b515a5f4c7dc03b38f27a9d60a49c8a3e1a1b91
size 3548
