version https://git-lfs.github.com/spec/v1
oid sha256:4210f177102cb6a4c29e51f54f5adf1dab153e6daf5797d4221244e5e32bdf49
size 6102
