version https://git-lfs.github.com/spec/v1
oid sha256:b4d5b3bb7cf97b5b36f83c6b12108177bb0bc61637223ea51811b38faae4d003
size 2778
